code_group_struct_t spec_decode_neg_8b10b_table_aa[code_group_t] = '{
	 // Negative CRD 
	10'b001111_0100  :  '{ 10'b001111_0100 ,  8'h1C , "K28_0" } , 
	10'b001111_1001  :  '{ 10'b001111_1001 ,  8'h3C , "K28_1" } , 
	10'b001111_0101  :  '{ 10'b001111_0101 ,  8'h5C , "K28_2" } , 
	10'b001111_0011  :  '{ 10'b001111_0011 ,  8'h7C , "K28_3" } , 
	10'b001111_0010  :  '{ 10'b001111_0010 ,  8'h9C , "K28_4" } , 
	10'b001111_1010  :  '{ 10'b001111_1010 ,  8'hBC , "K28_5" } , 
	10'b001111_0110  :  '{ 10'b001111_0110 ,  8'hDC , "K28_6" } , 
	10'b001111_1000  :  '{ 10'b001111_1000 ,  8'hFC , "K28_7" } , 
	10'b111010_1000  :  '{ 10'b111010_1000 ,  8'hF7 , "K23_7" } , 
	10'b110110_1000  :  '{ 10'b110110_1000 ,  8'hFB , "K27_7" } , 
	10'b101110_1000  :  '{ 10'b101110_1000 ,  8'hFD , "K29_7" } , 
	10'b011110_1000  :  '{ 10'b011110_1000 ,  8'hFE , "K30_7" }   
};


code_group_struct_t spec_decode_pos_8b10b_table_aa[code_group_t] = '{
	 // Positive CRD 
	10'b110000_1011  :  '{ 10'b110000_1011 ,  8'h1C , "K28_0" } , 
	10'b110000_0110  :  '{ 10'b110000_0110 ,  8'h3C , "K28_1" } , 
	10'b110000_1010  :  '{ 10'b110000_1010 ,  8'h5C , "K28_2" } , 
	10'b110000_1100  :  '{ 10'b110000_1100 ,  8'h7C , "K28_3" } , 
	10'b110000_1101  :  '{ 10'b110000_1101 ,  8'h9C , "K28_4" } , 
	10'b110000_0101  :  '{ 10'b110000_0101 ,  8'hBC , "K28_5" } , 
	10'b110000_1001  :  '{ 10'b110000_1001 ,  8'hDC , "K28_6" } , 
	10'b110000_0111  :  '{ 10'b110000_0111 ,  8'hFC , "K28_7" } , 
	10'b000101_0111  :  '{ 10'b000101_0111 ,  8'hF7 , "K23_7" } , 
	10'b001001_0111  :  '{ 10'b001001_0111 ,  8'hFB , "K27_7" } , 
	10'b010001_0111  :  '{ 10'b010001_0111 ,  8'hFD , "K29_7" } , 
	10'b100001_0111  :  '{ 10'b100001_0111 ,  8'hFE , "K30_7" }   
};


decode_table_t spec_decode_8b10b_table_aa[crd_t] = '{
	 NEGATIVE : spec_decode_neg_8b10b_table_aa,
	 POSITIVE : spec_decode_pos_8b10b_table_aa 
};


