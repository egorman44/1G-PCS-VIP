octet_t data_decode_neg_8b10b_table_aa[cg_t] = '{
	 // Negative CRD 
	10'b100111_0100  :   8'h00,  // "D0_0"
	10'b011101_0100  :   8'h01,  // "D1_0"
	10'b101101_0100  :   8'h02,  // "D2_0"
	10'b110001_1011  :   8'h03,  // "D3_0"
	10'b110101_0100  :   8'h04,  // "D4_0"
	10'b101001_1011  :   8'h05,  // "D5_0"
	10'b011001_1011  :   8'h06,  // "D6_0"
	10'b111000_1011  :   8'h07,  // "D7_0"
	10'b111001_0100  :   8'h08,  // "D8_0"
	10'b100101_1011  :   8'h09,  // "D9_0"
	10'b010101_1011  :   8'h0A,  // "D10_0"
	10'b110100_1011  :   8'h0B,  // "D11_0"
	10'b001101_1011  :   8'h0C,  // "D12_0"
	10'b101100_1011  :   8'h0D,  // "D13_0"
	10'b011100_1011  :   8'h0E,  // "D14_0"
	10'b010111_0100  :   8'h0F,  // "D15_0"
	10'b011011_0100  :   8'h10,  // "D16_0"
	10'b100011_1011  :   8'h11,  // "D17_0"
	10'b010011_1011  :   8'h12,  // "D18_0"
	10'b110010_1011  :   8'h13,  // "D19_0"
	10'b001011_1011  :   8'h14,  // "D20_0"
	10'b101010_1011  :   8'h15,  // "D21_0"
	10'b011010_1011  :   8'h16,  // "D22_0"
	10'b111010_0100  :   8'h17,  // "D23_0"
	10'b110011_0100  :   8'h18,  // "D24_0"
	10'b100110_1011  :   8'h19,  // "D25_0"
	10'b010110_1011  :   8'h1A,  // "D26_0"
	10'b110110_0100  :   8'h1B,  // "D27_0"
	10'b001110_1011  :   8'h1C,  // "D28_0"
	10'b101110_0100  :   8'h1D,  // "D29_0"
	10'b011110_0100  :   8'h1E,  // "D30_0"
	10'b101011_0100  :   8'h1F,  // "D31_0"
	10'b100111_1001  :   8'h20,  // "D0_1"
	10'b011101_1001  :   8'h21,  // "D1_1"
	10'b101101_1001  :   8'h22,  // "D2_1"
	10'b110001_1001  :   8'h23,  // "D3_1"
	10'b110101_1001  :   8'h24,  // "D4_1"
	10'b101001_1001  :   8'h25,  // "D5_1"
	10'b011001_1001  :   8'h26,  // "D6_1"
	10'b111000_1001  :   8'h27,  // "D7_1"
	10'b111001_1001  :   8'h28,  // "D8_1"
	10'b100101_1001  :   8'h29,  // "D9_1"
	10'b010101_1001  :   8'h2A,  // "D10_1"
	10'b110100_1001  :   8'h2B,  // "D11_1"
	10'b001101_1001  :   8'h2C,  // "D12_1"
	10'b101100_1001  :   8'h2D,  // "D13_1"
	10'b011100_1001  :   8'h2E,  // "D14_1"
	10'b010111_1001  :   8'h2F,  // "D15_1"
	10'b011011_1001  :   8'h30,  // "D16_1"
	10'b100011_1001  :   8'h31,  // "D17_1"
	10'b010011_1001  :   8'h32,  // "D18_1"
	10'b110010_1001  :   8'h33,  // "D19_1"
	10'b001011_1001  :   8'h34,  // "D20_1"
	10'b101010_1001  :   8'h35,  // "D21_1"
	10'b011010_1001  :   8'h36,  // "D22_1"
	10'b111010_1001  :   8'h37,  // "D23_1"
	10'b110011_1001  :   8'h38,  // "D24_1"
	10'b100110_1001  :   8'h39,  // "D25_1"
	10'b010110_1001  :   8'h3A,  // "D26_1"
	10'b110110_1001  :   8'h3B,  // "D27_1"
	10'b001110_1001  :   8'h3C,  // "D28_1"
	10'b101110_1001  :   8'h3D,  // "D29_1"
	10'b011110_1001  :   8'h3E,  // "D30_1"
	10'b101011_1001  :   8'h3F,  // "D31_1"
	10'b100111_0101  :   8'h40,  // "D0_2"
	10'b011101_0101  :   8'h41,  // "D1_2"
	10'b101101_0101  :   8'h42,  // "D2_2"
	10'b110001_0101  :   8'h43,  // "D3_2"
	10'b110101_0101  :   8'h44,  // "D4_2"
	10'b101001_0101  :   8'h45,  // "D5_2"
	10'b011001_0101  :   8'h46,  // "D6_2"
	10'b111000_0101  :   8'h47,  // "D7_2"
	10'b111001_0101  :   8'h48,  // "D8_2"
	10'b100101_0101  :   8'h49,  // "D9_2"
	10'b010101_0101  :   8'h4A,  // "D10_2"
	10'b110100_0101  :   8'h4B,  // "D11_2"
	10'b001101_0101  :   8'h4C,  // "D12_2"
	10'b101100_0101  :   8'h4D,  // "D13_2"
	10'b011100_0101  :   8'h4E,  // "D14_2"
	10'b010111_0101  :   8'h4F,  // "D15_2"
	10'b011011_0101  :   8'h50,  // "D16_2"
	10'b100011_0101  :   8'h51,  // "D17_2"
	10'b010011_0101  :   8'h52,  // "D18_2"
	10'b110010_0101  :   8'h53,  // "D19_2"
	10'b001011_0101  :   8'h54,  // "D20_2"
	10'b101010_0101  :   8'h55,  // "D21_2"
	10'b011010_0101  :   8'h56,  // "D22_2"
	10'b111010_0101  :   8'h57,  // "D23_2"
	10'b110011_0101  :   8'h58,  // "D24_2"
	10'b100110_0101  :   8'h59,  // "D25_2"
	10'b010110_0101  :   8'h5A,  // "D26_2"
	10'b110110_0101  :   8'h5B,  // "D27_2"
	10'b001110_0101  :   8'h5C,  // "D28_2"
	10'b101110_0101  :   8'h5D,  // "D29_2"
	10'b011110_0101  :   8'h5E,  // "D30_2"
	10'b101011_0101  :   8'h5F,  // "D31_2"
	10'b100111_0011  :   8'h60,  // "D0_3"
	10'b011101_0011  :   8'h61,  // "D1_3"
	10'b101101_0011  :   8'h62,  // "D2_3"
	10'b110001_1100  :   8'h63,  // "D3_3"
	10'b110101_0011  :   8'h64,  // "D4_3"
	10'b101001_1100  :   8'h65,  // "D5_3"
	10'b011001_1100  :   8'h66,  // "D6_3"
	10'b111000_1100  :   8'h67,  // "D7_3"
	10'b111001_0011  :   8'h68,  // "D8_3"
	10'b100101_1100  :   8'h69,  // "D9_3"
	10'b010101_1100  :   8'h6A,  // "D10_3"
	10'b110100_1100  :   8'h6B,  // "D11_3"
	10'b001101_1100  :   8'h6C,  // "D12_3"
	10'b101100_1100  :   8'h6D,  // "D13_3"
	10'b011100_1100  :   8'h6E,  // "D14_3"
	10'b010111_0011  :   8'h6F,  // "D15_3"
	10'b011011_0011  :   8'h70,  // "D16_3"
	10'b100011_1100  :   8'h71,  // "D17_3"
	10'b010011_1100  :   8'h72,  // "D18_3"
	10'b110010_1100  :   8'h73,  // "D19_3"
	10'b001011_1100  :   8'h74,  // "D20_3"
	10'b101010_1100  :   8'h75,  // "D21_3"
	10'b011010_1100  :   8'h76,  // "D22_3"
	10'b111010_0011  :   8'h77,  // "D23_3"
	10'b110011_0011  :   8'h78,  // "D24_3"
	10'b100110_1100  :   8'h79,  // "D25_3"
	10'b010110_1100  :   8'h7A,  // "D26_3"
	10'b110110_0011  :   8'h7B,  // "D27_3"
	10'b001110_1100  :   8'h7C,  // "D28_3"
	10'b101110_0011  :   8'h7D,  // "D29_3"
	10'b011110_0011  :   8'h7E,  // "D30_3"
	10'b101011_0011  :   8'h7F,  // "D31_3"
	10'b100111_0010  :   8'h80,  // "D0_4"
	10'b011101_0010  :   8'h81,  // "D1_4"
	10'b101101_0010  :   8'h82,  // "D2_4"
	10'b110001_1101  :   8'h83,  // "D3_4"
	10'b110101_0010  :   8'h84,  // "D4_4"
	10'b101001_1101  :   8'h85,  // "D5_4" 1000_0101
	10'b011001_1101  :   8'h86,  // "D6_4"
	10'b111000_1101  :   8'h87,  // "D7_4"
	10'b111001_0010  :   8'h88,  // "D8_4"
	10'b100101_1101  :   8'h89,  // "D9_4"
	10'b010101_1101  :   8'h8A,  // "D10_4"
	10'b110100_1101  :   8'h8B,  // "D11_4"
	10'b001101_1101  :   8'h8C,  // "D12_4"
	10'b101100_1101  :   8'h8D,  // "D13_4"
	10'b011100_1101  :   8'h8E,  // "D14_4"
	10'b010111_0010  :   8'h8F,  // "D15_4"
	10'b011011_0010  :   8'h90,  // "D16_4"
	10'b100011_1101  :   8'h91,  // "D17_4"
	10'b010011_1101  :   8'h92,  // "D18_4"
	10'b110010_1101  :   8'h93,  // "D19_4"
	10'b001011_1101  :   8'h94,  // "D20_4"
	10'b101010_1101  :   8'h95,  // "D21_4"
	10'b011010_1101  :   8'h96,  // "D22_4"
	10'b111010_0010  :   8'h97,  // "D23_4"
	10'b110011_0010  :   8'h98,  // "D24_4"
	10'b100110_1101  :   8'h99,  // "D25_4"
	10'b010110_1101  :   8'h9A,  // "D26_4"
	10'b110110_0010  :   8'h9B,  // "D27_4"
	10'b001110_1101  :   8'h9C,  // "D28_4"
	10'b101110_0010  :   8'h9D,  // "D29_4"
	10'b011110_0010  :   8'h9E,  // "D30_4"
	10'b101011_0010  :   8'h9F,  // "D31_4"
	10'b100111_1010  :   8'hA0,  // "D0_5"
	10'b011101_1010  :   8'hA1,  // "D1_5"
	10'b101101_1010  :   8'hA2,  // "D2_5"
	10'b110001_1010  :   8'hA3,  // "D3_5"
	10'b110101_1010  :   8'hA4,  // "D4_5"
	10'b101001_1010  :   8'hA5,  // "D5_5"
	10'b011001_1010  :   8'hA6,  // "D6_5"
	10'b111000_1010  :   8'hA7,  // "D7_5"
	10'b111001_1010  :   8'hA8,  // "D8_5"
	10'b100101_1010  :   8'hA9,  // "D9_5"
	10'b010101_1010  :   8'hAA,  // "D10_5"
	10'b110100_1010  :   8'hAB,  // "D11_5"
	10'b001101_1010  :   8'hAC,  // "D12_5"
	10'b101100_1010  :   8'hAD,  // "D13_5"
	10'b011100_1010  :   8'hAE,  // "D14_5"
	10'b010111_1010  :   8'hAF,  // "D15_5"
	10'b011011_1010  :   8'hB0,  // "D16_5"
	10'b100011_1010  :   8'hB1,  // "D17_5"
	10'b010011_1010  :   8'hB2,  // "D18_5"
	10'b110010_1010  :   8'hB3,  // "D19_5"
	10'b001011_1010  :   8'hB4,  // "D20_5"
	10'b101010_1010  :   8'hB5,  // "D21_5"
	10'b011010_1010  :   8'hB6,  // "D22_5"
	10'b111010_1010  :   8'hB7,  // "D23_5"
	10'b110011_1010  :   8'hB8,  // "D24_5"
	10'b100110_1010  :   8'hB9,  // "D25_5"
	10'b010110_1010  :   8'hBA,  // "D26_5"
	10'b110110_1010  :   8'hBB,  // "D27_5"
	10'b001110_1010  :   8'hBC,  // "D28_5"
	10'b101110_1010  :   8'hBD,  // "D29_5"
	10'b011110_1010  :   8'hBE,  // "D30_5"
	10'b101011_1010  :   8'hBF,  // "D31_5"
	10'b100111_0110  :   8'hC0,  // "D0_6"
	10'b011101_0110  :   8'hC1,  // "D1_6"
	10'b101101_0110  :   8'hC2,  // "D2_6"
	10'b110001_0110  :   8'hC3,  // "D3_6"
	10'b110101_0110  :   8'hC4,  // "D4_6"
	10'b101001_0110  :   8'hC5,  // "D5_6"
	10'b011001_0110  :   8'hC6,  // "D6_6"
	10'b111000_0110  :   8'hC7,  // "D7_6"
	10'b111001_0110  :   8'hC8,  // "D8_6"
	10'b100101_0110  :   8'hC9,  // "D9_6"
	10'b010101_0110  :   8'hCA,  // "D10_6"
	10'b110100_0110  :   8'hCB,  // "D11_6"
	10'b001101_0110  :   8'hCC,  // "D12_6"
	10'b101100_0110  :   8'hCD,  // "D13_6"
	10'b011100_0110  :   8'hCE,  // "D14_6"
	10'b010111_0110  :   8'hCF,  // "D15_6"
	10'b011011_0110  :   8'hD0,  // "D16_6"
	10'b100011_0110  :   8'hD1,  // "D17_6"
	10'b010011_0110  :   8'hD2,  // "D18_6"
	10'b110010_0110  :   8'hD3,  // "D19_6"
	10'b001011_0110  :   8'hD4,  // "D20_6"
	10'b101010_0110  :   8'hD5,  // "D21_6"
	10'b011010_0110  :   8'hD6,  // "D22_6"
	10'b111010_0110  :   8'hD7,  // "D23_6"
	10'b110011_0110  :   8'hD8,  // "D24_6"
	10'b100110_0110  :   8'hD9,  // "D25_6"
	10'b010110_0110  :   8'hDA,  // "D26_6"
	10'b110110_0110  :   8'hDB,  // "D27_6"
	10'b001110_0110  :   8'hDC,  // "D28_6"
	10'b101110_0110  :   8'hDD,  // "D29_6"
	10'b011110_0110  :   8'hDE,  // "D30_6"
	10'b101011_0110  :   8'hDF,  // "D31_6"
	10'b100111_0001  :   8'hE0,  // "D0_7"
	10'b011101_0001  :   8'hE1,  // "D1_7"
	10'b101101_0001  :   8'hE2,  // "D2_7"
	10'b110001_1110  :   8'hE3,  // "D3_7"
	10'b110101_0001  :   8'hE4,  // "D4_7"
	10'b101001_1110  :   8'hE5,  // "D5_7"
	10'b011001_1110  :   8'hE6,  // "D6_7"
	10'b111000_1110  :   8'hE7,  // "D7_7"
	10'b111001_0001  :   8'hE8,  // "D8_7"
	10'b100101_1110  :   8'hE9,  // "D9_7"
	10'b010101_1110  :   8'hEA,  // "D10_7"
	10'b110100_1110  :   8'hEB,  // "D11_7"
	10'b001101_1110  :   8'hEC,  // "D12_7"
	10'b101100_1110  :   8'hED,  // "D13_7"
	10'b011100_1110  :   8'hEE,  // "D14_7"
	10'b010111_0001  :   8'hEF,  // "D15_7"
	10'b011011_0001  :   8'hF0,  // "D16_7"
	10'b100011_0111  :   8'hF1,  // "D17_7"
	10'b010011_0111  :   8'hF2,  // "D18_7"
	10'b110010_1110  :   8'hF3,  // "D19_7"
	10'b001011_0111  :   8'hF4,  // "D20_7"
	10'b101010_1110  :   8'hF5,  // "D21_7"
	10'b011010_1110  :   8'hF6,  // "D22_7"
	10'b111010_0001  :   8'hF7,  // "D23_7"
	10'b110011_0001  :   8'hF8,  // "D24_7"
	10'b100110_1110  :   8'hF9,  // "D25_7"
	10'b010110_1110  :   8'hFA,  // "D26_7"
	10'b110110_0001  :   8'hFB,  // "D27_7"
	10'b001110_1110  :   8'hFC,  // "D28_7"
	10'b101110_0001  :   8'hFD,  // "D29_7"
	10'b011110_0001  :   8'hFE,  // "D30_7"
	10'b101011_0001  :   8'hFF   // "D31_7"
};


octet_t data_decode_pos_8b10b_table_aa[cg_t] = '{
	 // Positive CRD 
	10'b011000_1011  :   8'h00,  // "D0_0"
	10'b100010_1011  :   8'h01,  // "D1_0"
	10'b010010_1011  :   8'h02,  // "D2_0"
	10'b110001_0100  :   8'h03,  // "D3_0"
	10'b001010_1011  :   8'h04,  // "D4_0"
	10'b101001_0100  :   8'h05,  // "D5_0"
	10'b011001_0100  :   8'h06,  // "D6_0"
	10'b000111_0100  :   8'h07,  // "D7_0"
	10'b000110_1011  :   8'h08,  // "D8_0"
	10'b100101_0100  :   8'h09,  // "D9_0"
	10'b010101_0100  :   8'h0A,  // "D10_0"
	10'b110100_0100  :   8'h0B,  // "D11_0"
	10'b001101_0100  :   8'h0C,  // "D12_0"
	10'b101100_0100  :   8'h0D,  // "D13_0"
	10'b011100_0100  :   8'h0E,  // "D14_0"
	10'b101000_1011  :   8'h0F,  // "D15_0"
	10'b100100_1011  :   8'h10,  // "D16_0"
	10'b100011_0100  :   8'h11,  // "D17_0"
	10'b010011_0100  :   8'h12,  // "D18_0"
	10'b110010_0100  :   8'h13,  // "D19_0"
	10'b001011_0100  :   8'h14,  // "D20_0"
	10'b101010_0100  :   8'h15,  // "D21_0"
	10'b011010_0100  :   8'h16,  // "D22_0"
	10'b000101_1011  :   8'h17,  // "D23_0"
	10'b001100_1011  :   8'h18,  // "D24_0"
	10'b100110_0100  :   8'h19,  // "D25_0"
	10'b010110_0100  :   8'h1A,  // "D26_0"
	10'b001001_1011  :   8'h1B,  // "D27_0"
	10'b001110_0100  :   8'h1C,  // "D28_0"
	10'b010001_1011  :   8'h1D,  // "D29_0"
	10'b100001_1011  :   8'h1E,  // "D30_0"
	10'b010100_1011  :   8'h1F,  // "D31_0"
	10'b011000_1001  :   8'h20,  // "D0_1"
	10'b100010_1001  :   8'h21,  // "D1_1"
	10'b010010_1001  :   8'h22,  // "D2_1"
	10'b110001_1001  :   8'h23,  // "D3_1"
	10'b001010_1001  :   8'h24,  // "D4_1"
	10'b101001_1001  :   8'h25,  // "D5_1"
	10'b011001_1001  :   8'h26,  // "D6_1"
	10'b000111_1001  :   8'h27,  // "D7_1"
	10'b000110_1001  :   8'h28,  // "D8_1"
	10'b100101_1001  :   8'h29,  // "D9_1"
	10'b010101_1001  :   8'h2A,  // "D10_1"
	10'b110100_1001  :   8'h2B,  // "D11_1"
	10'b001101_1001  :   8'h2C,  // "D12_1"
	10'b101100_1001  :   8'h2D,  // "D13_1"
	10'b011100_1001  :   8'h2E,  // "D14_1"
	10'b101000_1001  :   8'h2F,  // "D15_1"
	10'b100100_1001  :   8'h30,  // "D16_1"
	10'b100011_1001  :   8'h31,  // "D17_1"
	10'b010011_1001  :   8'h32,  // "D18_1"
	10'b110010_1001  :   8'h33,  // "D19_1"
	10'b001011_1001  :   8'h34,  // "D20_1"
	10'b101010_1001  :   8'h35,  // "D21_1"
	10'b011010_1001  :   8'h36,  // "D22_1"
	10'b000101_1001  :   8'h37,  // "D23_1"
	10'b001100_1001  :   8'h38,  // "D24_1"
	10'b100110_1001  :   8'h39,  // "D25_1"
	10'b010110_1001  :   8'h3A,  // "D26_1"
	10'b001001_1001  :   8'h3B,  // "D27_1"
	10'b001110_1001  :   8'h3C,  // "D28_1"
	10'b010001_1001  :   8'h3D,  // "D29_1"
	10'b100001_1001  :   8'h3E,  // "D30_1"
	10'b010100_1001  :   8'h3F,  // "D31_1"
	10'b011000_0101  :   8'h40,  // "D0_2"
	10'b100010_0101  :   8'h41,  // "D1_2"
	10'b010010_0101  :   8'h42,  // "D2_2"
	10'b110001_0101  :   8'h43,  // "D3_2"
	10'b001010_0101  :   8'h44,  // "D4_2"
	10'b101001_0101  :   8'h45,  // "D5_2"
	10'b011001_0101  :   8'h46,  // "D6_2"
	10'b000111_0101  :   8'h47,  // "D7_2"
	10'b000110_0101  :   8'h48,  // "D8_2"
	10'b100101_0101  :   8'h49,  // "D9_2"
	10'b010101_0101  :   8'h4A,  // "D10_2"
	10'b110100_0101  :   8'h4B,  // "D11_2"
	10'b001101_0101  :   8'h4C,  // "D12_2"
	10'b101100_0101  :   8'h4D,  // "D13_2"
	10'b011100_0101  :   8'h4E,  // "D14_2"
	10'b101000_0101  :   8'h4F,  // "D15_2"
	10'b100100_0101  :   8'h50,  // "D16_2"
	10'b100011_0101  :   8'h51,  // "D17_2"
	10'b010011_0101  :   8'h52,  // "D18_2"
	10'b110010_0101  :   8'h53,  // "D19_2"
	10'b001011_0101  :   8'h54,  // "D20_2"
	10'b101010_0101  :   8'h55,  // "D21_2"
	10'b011010_0101  :   8'h56,  // "D22_2"
	10'b000101_0101  :   8'h57,  // "D23_2"
	10'b001100_0101  :   8'h58,  // "D24_2"
	10'b100110_0101  :   8'h59,  // "D25_2"
	10'b010110_0101  :   8'h5A,  // "D26_2"
	10'b001001_0101  :   8'h5B,  // "D27_2"
	10'b001110_0101  :   8'h5C,  // "D28_2"
	10'b010001_0101  :   8'h5D,  // "D29_2"
	10'b100001_0101  :   8'h5E,  // "D30_2"
	10'b010100_0101  :   8'h5F,  // "D31_2"
	10'b011000_1100  :   8'h60,  // "D0_3"
	10'b100010_1100  :   8'h61,  // "D1_3"
	10'b010010_1100  :   8'h62,  // "D2_3"
	10'b110001_0011  :   8'h63,  // "D3_3"
	10'b001010_1100  :   8'h64,  // "D4_3"
	10'b101001_0011  :   8'h65,  // "D5_3"
	10'b011001_0011  :   8'h66,  // "D6_3"
	10'b000111_0011  :   8'h67,  // "D7_3"
	10'b000110_1100  :   8'h68,  // "D8_3"
	10'b100101_0011  :   8'h69,  // "D9_3"
	10'b010101_0011  :   8'h6A,  // "D10_3"
	10'b110100_0011  :   8'h6B,  // "D11_3"
	10'b001101_0011  :   8'h6C,  // "D12_3"
	10'b101100_0011  :   8'h6D,  // "D13_3"
	10'b011100_0011  :   8'h6E,  // "D14_3"
	10'b101000_1100  :   8'h6F,  // "D15_3"
	10'b100100_1100  :   8'h70,  // "D16_3"
	10'b100011_0011  :   8'h71,  // "D17_3"
	10'b010011_0011  :   8'h72,  // "D18_3"
	10'b110010_0011  :   8'h73,  // "D19_3"
	10'b001011_0011  :   8'h74,  // "D20_3"
	10'b101010_0011  :   8'h75,  // "D21_3"
	10'b011010_0011  :   8'h76,  // "D22_3"
	10'b000101_1100  :   8'h77,  // "D23_3"
	10'b001100_1100  :   8'h78,  // "D24_3"
	10'b100110_0011  :   8'h79,  // "D25_3"
	10'b010110_0011  :   8'h7A,  // "D26_3"
	10'b001001_1100  :   8'h7B,  // "D27_3"
	10'b001110_0011  :   8'h7C,  // "D28_3"
	10'b010001_1100  :   8'h7D,  // "D29_3"
	10'b100001_1100  :   8'h7E,  // "D30_3"
	10'b010100_1100  :   8'h7F,  // "D31_3"
	10'b011000_1101  :   8'h80,  // "D0_4"
	10'b100010_1101  :   8'h81,  // "D1_4"
	10'b010010_1101  :   8'h82,  // "D2_4"
	10'b110001_0010  :   8'h83,  // "D3_4"
	10'b001010_1101  :   8'h84,  // "D4_4"
	10'b101001_0010  :   8'h85,  // "D5_4"
	10'b011001_0010  :   8'h86,  // "D6_4"
	10'b000111_0010  :   8'h87,  // "D7_4"
	10'b000110_1101  :   8'h88,  // "D8_4"
	10'b100101_0010  :   8'h89,  // "D9_4"
	10'b010101_0010  :   8'h8A,  // "D10_4"
	10'b110100_0010  :   8'h8B,  // "D11_4"
	10'b001101_0010  :   8'h8C,  // "D12_4"
	10'b101100_0010  :   8'h8D,  // "D13_4"
	10'b011100_0010  :   8'h8E,  // "D14_4"
	10'b101000_1101  :   8'h8F,  // "D15_4"
	10'b100100_1101  :   8'h90,  // "D16_4"
	10'b100011_0010  :   8'h91,  // "D17_4"
	10'b010011_0010  :   8'h92,  // "D18_4"
	10'b110010_0010  :   8'h93,  // "D19_4"
	10'b001011_0010  :   8'h94,  // "D20_4"
	10'b101010_0010  :   8'h95,  // "D21_4"
	10'b011010_0010  :   8'h96,  // "D22_4"
	10'b000101_1101  :   8'h97,  // "D23_4"
	10'b001100_1101  :   8'h98,  // "D24_4"
	10'b100110_0010  :   8'h99,  // "D25_4"
	10'b010110_0010  :   8'h9A,  // "D26_4"
	10'b001001_1101  :   8'h9B,  // "D27_4"
	10'b001110_0010  :   8'h9C,  // "D28_4"
	10'b010001_1101  :   8'h9D,  // "D29_4"
	10'b100001_1101  :   8'h9E,  // "D30_4"
	10'b010100_1101  :   8'h9F,  // "D31_4"
	10'b011000_1010  :   8'hA0,  // "D0_5"
	10'b100010_1010  :   8'hA1,  // "D1_5"
	10'b010010_1010  :   8'hA2,  // "D2_5"
	10'b110001_1010  :   8'hA3,  // "D3_5"
	10'b001010_1010  :   8'hA4,  // "D4_5"
	10'b101001_1010  :   8'hA5,  // "D5_5"
	10'b011001_1010  :   8'hA6,  // "D6_5"
	10'b000111_1010  :   8'hA7,  // "D7_5"
	10'b000110_1010  :   8'hA8,  // "D8_5"
	10'b100101_1010  :   8'hA9,  // "D9_5"
	10'b010101_1010  :   8'hAA,  // "D10_5"
	10'b110100_1010  :   8'hAB,  // "D11_5"
	10'b001101_1010  :   8'hAC,  // "D12_5"
	10'b101100_1010  :   8'hAD,  // "D13_5"
	10'b011100_1010  :   8'hAE,  // "D14_5"
	10'b101000_1010  :   8'hAF,  // "D15_5"
	10'b100100_1010  :   8'hB0,  // "D16_5"
	10'b100011_1010  :   8'hB1,  // "D17_5"
	10'b010011_1010  :   8'hB2,  // "D18_5"
	10'b110010_1010  :   8'hB3,  // "D19_5"
	10'b001011_1010  :   8'hB4,  // "D20_5"
	10'b101010_1010  :   8'hB5,  // "D21_5"
	10'b011010_1010  :   8'hB6,  // "D22_5"
	10'b000101_1010  :   8'hB7,  // "D23_5"
	10'b001100_1010  :   8'hB8,  // "D24_5"
	10'b100110_1010  :   8'hB9,  // "D25_5"
	10'b010110_1010  :   8'hBA,  // "D26_5"
	10'b001001_1010  :   8'hBB,  // "D27_5"
	10'b001110_1010  :   8'hBC,  // "D28_5"
	10'b010001_1010  :   8'hBD,  // "D29_5"
	10'b100001_1010  :   8'hBE,  // "D30_5"
	10'b010100_1010  :   8'hBF,  // "D31_5"
	10'b011000_0110  :   8'hC0,  // "D0_6"
	10'b100010_0110  :   8'hC1,  // "D1_6"
	10'b010010_0110  :   8'hC2,  // "D2_6"
	10'b110001_0110  :   8'hC3,  // "D3_6"
	10'b001010_0110  :   8'hC4,  // "D4_6"
	10'b101001_0110  :   8'hC5,  // "D5_6"
	10'b011001_0110  :   8'hC6,  // "D6_6"
	10'b000111_0110  :   8'hC7,  // "D7_6"
	10'b000110_0110  :   8'hC8,  // "D8_6"
	10'b100101_0110  :   8'hC9,  // "D9_6"
	10'b010101_0110  :   8'hCA,  // "D10_6"
	10'b110100_0110  :   8'hCB,  // "D11_6"
	10'b001101_0110  :   8'hCC,  // "D12_6"
	10'b101100_0110  :   8'hCD,  // "D13_6"
	10'b011100_0110  :   8'hCE,  // "D14_6"
	10'b101000_0110  :   8'hCF,  // "D15_6"
	10'b100100_0110  :   8'hD0,  // "D16_6"
	10'b100011_0110  :   8'hD1,  // "D17_6"
	10'b010011_0110  :   8'hD2,  // "D18_6"
	10'b110010_0110  :   8'hD3,  // "D19_6"
	10'b001011_0110  :   8'hD4,  // "D20_6"
	10'b101010_0110  :   8'hD5,  // "D21_6"
	10'b011010_0110  :   8'hD6,  // "D22_6"
	10'b000101_0110  :   8'hD7,  // "D23_6"
	10'b001100_0110  :   8'hD8,  // "D24_6"
	10'b100110_0110  :   8'hD9,  // "D25_6"
	10'b010110_0110  :   8'hDA,  // "D26_6"
	10'b001001_0110  :   8'hDB,  // "D27_6"
	10'b001110_0110  :   8'hDC,  // "D28_6"
	10'b010001_0110  :   8'hDD,  // "D29_6"
	10'b100001_0110  :   8'hDE,  // "D30_6"
	10'b010100_0110  :   8'hDF,  // "D31_6"
	10'b011000_1110  :   8'hE0,  // "D0_7"
	10'b100010_1110  :   8'hE1,  // "D1_7"
	10'b010010_1110  :   8'hE2,  // "D2_7"
	10'b110001_0001  :   8'hE3,  // "D3_7"
	10'b001010_1110  :   8'hE4,  // "D4_7"
	10'b101001_0001  :   8'hE5,  // "D5_7"
	10'b011001_0001  :   8'hE6,  // "D6_7"
	10'b000111_0001  :   8'hE7,  // "D7_7"
	10'b000110_1110  :   8'hE8,  // "D8_7"
	10'b100101_0001  :   8'hE9,  // "D9_7"
	10'b010101_0001  :   8'hEA,  // "D10_7"
	10'b110100_1000  :   8'hEB,  // "D11_7"
	10'b001101_0001  :   8'hEC,  // "D12_7"
	10'b101100_1000  :   8'hED,  // "D13_7"
	10'b011100_1000  :   8'hEE,  // "D14_7"
	10'b101000_1110  :   8'hEF,  // "D15_7"
	10'b100100_1110  :   8'hF0,  // "D16_7"
	10'b100011_0001  :   8'hF1,  // "D17_7"
	10'b010011_0001  :   8'hF2,  // "D18_7"
	10'b110010_0001  :   8'hF3,  // "D19_7"
	10'b001011_0001  :   8'hF4,  // "D20_7"
	10'b101010_0001  :   8'hF5,  // "D21_7"
	10'b011010_0001  :   8'hF6,  // "D22_7"
	10'b000101_1110  :   8'hF7,  // "D23_7"
	10'b001100_1110  :   8'hF8,  // "D24_7"
	10'b100110_0001  :   8'hF9,  // "D25_7"
	10'b010110_0001  :   8'hFA,  // "D26_7"
	10'b001001_1110  :   8'hFB,  // "D27_7"
	10'b001110_0001  :   8'hFC,  // "D28_7"
	10'b010001_1110  :   8'hFD,  // "D29_7"
	10'b100001_1110  :   8'hFE,  // "D30_7"
	10'b010100_1110  :   8'hFF   // "D31_7"
};


decode_table_t data_decode_8b10b_table_aa[crd_t] = '{
	 NEGATIVE : data_decode_neg_8b10b_table_aa,
	 POSITIVE : data_decode_pos_8b10b_table_aa 
};


octet_t spec_decode_neg_8b10b_table_aa[cg_t] = '{
	 // Negative CRD 
	10'b001111_0100  :   8'h1C,  // "K28_0"
	10'b001111_1001  :   8'h3C,  // "K28_1"
	10'b001111_0101  :   8'h5C,  // "K28_2"
	10'b001111_0011  :   8'h7C,  // "K28_3"
	10'b001111_0010  :   8'h9C,  // "K28_4"
	10'b001111_1010  :   8'hBC,  // "K28_5"
	10'b001111_0110  :   8'hDC,  // "K28_6"
	10'b001111_1000  :   8'hFC,  // "K28_7"
	10'b111010_1000  :   8'hF7,  // "K23_7"
	10'b110110_1000  :   8'hFB,  // "K27_7"
	10'b101110_1000  :   8'hFD,  // "K29_7"
	10'b011110_1000  :   8'hFE   // "K30_7"
};


octet_t spec_decode_pos_8b10b_table_aa[cg_t] = '{
	 // Positive CRD 
	10'b110000_1011  :   8'h1C,  // "K28_0"
	10'b110000_0110  :   8'h3C,  // "K28_1"
	10'b110000_1010  :   8'h5C,  // "K28_2"
	10'b110000_1100  :   8'h7C,  // "K28_3"
	10'b110000_1101  :   8'h9C,  // "K28_4"
	10'b110000_0101  :   8'hBC,  // "K28_5"
	10'b110000_1001  :   8'hDC,  // "K28_6"
	10'b110000_0111  :   8'hFC,  // "K28_7"
	10'b000101_0111  :   8'hF7,  // "K23_7"
	10'b001001_0111  :   8'hFB,  // "K27_7"
	10'b010001_0111  :   8'hFD,  // "K29_7"
	10'b100001_0111  :   8'hFE   // "K30_7"
};


decode_table_t spec_decode_8b10b_table_aa[crd_t] = '{
	 NEGATIVE : spec_decode_neg_8b10b_table_aa,
	 POSITIVE : spec_decode_pos_8b10b_table_aa 
};


